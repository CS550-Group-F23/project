`include "def.vh"
module array_top (
    input clk,
    input [`DW-1:0] A [`SZ*`SZ-1:0],
    input [`DW-1:0] W [`SZ-1:0],
    output [`DW-1:0] O,
    input ready,
    output valid
);


    
endmodule