`define DW 16
`define SZ 3
`define SZ_D $clog2(`SZ)
`define BLOCK `SZ*`DW