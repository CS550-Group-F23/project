`define DW 16
`define SZ 3